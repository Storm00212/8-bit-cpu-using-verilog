// ============================================================================
// CPU Top-Level Module
// ============================================================================
// 
// The CPU Top-Level Module integrates all the individual components of the
// 8-bit CPU into a complete, functional processor. It provides the external
// interface and handles the interconnection between components.
// 
// Component Connections:
// - Control Unit orchestrates all operations
// - Register File stores CPU state
// - ALU performs calculations
// - RAM stores data
// - ROM stores program code
// 
// Bus Architecture:
// - 8-bit bidirectional data bus
// - 16-bit unidirectional address bus
// - Separate ROM and RAM address spaces
// ============================================================================

`include "instructions.vh"

module cpu_top (
    // External Interface
    input wire clk,           // System clock - all operations synchronous
    input wire reset,         // Asynchronous reset - initializes CPU
    
    // Bus Interface
    output wire [7:0] data_bus,      // 8-bit bidirectional data bus
    output wire [15:0] addr_bus,     // 16-bit address bus (output only)
    output wire mem_read,            // Memory read enable
    output wire mem_write,           // Memory write enable
    
    // Debug/Status Outputs
    output wire [7:0] acc_out,      // Accumulator value (debug)
    output wire [15:0] pc_out,      // Program counter value (debug)
    output wire [7:0] flags_out,     // Flags register (debug)
    output wire [7:0] x_out,         // X register value (debug)
    output wire [7:0] y_out,         // Y register value (debug)
    output wire halt                 // CPU halt status
);

    // =========================================================================
    // Signal Declarations
    // =========================================================================
    
    // -------------------- Control Signals --------------------
    // These signals are generated by the Control Unit and control
    // the operation of other CPU components.
    
    wire acc_write, x_write, y_write;      // Register write enables
    wire pc_write, pc_inc, pc_load;       // PC control signals
    wire sp_write, ir_write, flags_write;  // Register write enables
    wire alu_done;                          // ALU operation complete
    wire done;                              // Instruction complete
    wire [3:0] alu_operation;              // ALU operation code
    wire [15:0] pc_direct;                 // Direct PC value for jumps
    
    // -------------------- Data Signals --------------------
    // These signals carry data between CPU components.
    
    wire [7:0] acc_reg, x_reg, y_reg;      // Register values
    wire [7:0] sp_reg, ir_reg, flags_reg; // Register values
    wire [15:0] pc_reg;                   // Program counter
    reg [15:0] pc_current;               // Current PC value (registered)
    
    // -------------------- Memory Interface --------------------
    // These signals interface with ROM and RAM modules.
    
    wire [7:0] ram_data_out, rom_data_out; // Memory data outputs
    wire ram_ready;                         // RAM ready signal
    wire [15:0] mem_addr;                  // Memory address
    
    wire mem_data_from_ram;                 // Data source selection
    wire mem_data_from_rom;                 // Data source selection
    
    // -------------------- ALU Signals --------------------
    wire [7:0] alu_result;                 // ALU result output
    wire [7:0] alu_flags;                  // ALU flags output
    
    // =========================================================================
    // PC Register - Captures PC value for control unit
    // =========================================================================
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            pc_current <= 16'd0;
        end else begin
            pc_current <= pc_reg;
        end
    end
    
    // =========================================================================
    // Module Instantiations
    // =========================================================================
    
    // -------------------- Register File --------------------
    // The Register File stores all CPU registers including the accumulator,
    // index registers (X, Y), program counter, stack pointer, instruction
    // register, and flags register.
    //
    // Inputs:
    //   - clk, reset: Clock and reset signals
    //   - data_in: Data to write to registers
    //   - Various write enable signals
    //   - PC control signals
    //
    // Outputs:
    //   - acc_out, x_out, y_out, pc_out, sp_out, ir_out, flags_out
    //   - addr_bus: Address for memory operations
    
    register_file reg_file (
        .clk(clk),
        .reset(reset),
        .data_in(data_bus),
        .acc_write(acc_write),
        .x_write(x_write),
        .y_write(y_write),
        .pc_write(pc_write),
        .sp_write(sp_write),
        .ir_write(ir_write),
        .flags_write(flags_write),
        .pc_direct(pc_direct),
        .pc_inc(pc_inc),
        .pc_load(pc_load),
        .acc_out(acc_reg),
        .x_out(x_reg),
        .y_out(y_reg),
        .pc_out(pc_reg),
        .sp_out(sp_reg),
        .ir_out(ir_reg),
        .flags_out(flags_reg),
        .addr_bus(addr_bus)
    );
    
    // -------------------- ALU (Arithmetic Logic Unit) --------------------
    // The ALU performs all arithmetic, logical, and mathematical operations.
    // It receives operands from the register file and returns results and flags.
    //
    // Inputs:
    //   - a: First operand (typically accumulator)
    //   - b: Second operand (from data bus)
    //   - operation: Operation code
    //   - clk, reset: Clock and reset
    //
    // Outputs:
    //   - result: Operation result
    //   - flags: Status flags
    //   - done: Operation complete signal
    
    alu alu_unit (
        .clk(clk),
        .reset(reset),
        .a(acc_reg),
        .b(data_bus),
        .operation(alu_operation),
        .result(alu_result),
        .flags(alu_flags),
        .done(alu_done)
    );
    
    // -------------------- Control Unit --------------------
    // The Control Unit decodes instructions and generates control signals.
    // It orchestrates the operation of all other CPU components.
    //
    // Inputs:
    //   - clk, reset: Clock and reset
    //   - opcode: Current instruction opcode
    //   - flags_in: Current flags register value
    //   - alu_done: ALU operation complete
    //   - data_bus: Data from memory
    //   - pc_current: Current PC value
    //
    // Outputs:
    //   - Various control signals to other components
    //   - done: Instruction complete
    
    control_unit cu (
        .clk(clk),
        .reset(reset),
        .opcode(data_bus),
        .flags_in(flags_reg),
        .alu_done(alu_done),
        .data_bus(data_bus),
        .pc_current(pc_current),
        .alu_operation(alu_operation),
        .acc_write(acc_write),
        .x_write(x_write),
        .y_write(y_write),
        .pc_write(pc_write),
        .pc_inc(pc_inc),
        .pc_load(pc_load),
        .pc_direct(pc_direct),
        .sp_write(sp_write),
        .ir_write(ir_write),
        .flags_write(flags_write),
        .mem_read(mem_data_from_rom),
        .mem_write(mem_write),
        .mem_addr(mem_addr),
        .done(done)
    );
    
    // -------------------- RAM Module --------------------
    // Random Access Memory provides volatile data storage for the CPU.
    // All addresses except 0x0000-0x00FF access RAM.
    //
    // Inputs:
    //   - clk, reset: Clock and reset
    //   - addr: Memory address
    //   - data_in: Data to write
    //   - write_enable, read_enable: Control signals
    //
    // Outputs:
    //   - data_out: Data read from memory
    //   - ready: Memory ready signal
    
    ram ram_module (
        .clk(clk),
        .reset(reset),
        .addr(addr_bus),
        .data_in(acc_reg),
        .write_enable(mem_write),
        .read_enable(mem_data_from_ram),
        .data_out(ram_data_out),
        .ready(ram_ready)
    );
    
    // -------------------- ROM Module --------------------
    // Read-Only Memory stores the program code. Addresses 0x0000-0x00FF
    // access ROM for instruction fetch.
    //
    // Inputs:
    //   - addr: Memory address
    //
    // Outputs:
    //   - data_out: Instruction byte
    
    rom rom_module (
        .addr(addr_bus),
        .data_out(rom_data_out)
    );
    
    // =========================================================================
    // Memory Interface Logic
    // =========================================================================
    
    // -------------------- Memory Source Selection --------------------
    // The CPU uses a simple memory map to determine whether to access
    // ROM or RAM based on the address.
    //
    // Memory Map:
    //   0x0000 - 0x00FF: ROM (Program memory)
    //   0x0100 - 0xFFFF: RAM (Data memory)
    //
    // Note: This is a simplified design. A more complex design might
    // use memory-mapped I/O or have separate instruction and data caches.
    
    // ROM is accessed for addresses in the first 256 bytes
    assign mem_data_from_rom = (addr_bus[15:8] == 8'h00);
    
    // RAM is accessed for all other addresses
    assign mem_data_from_ram = (addr_bus[15:8] != 8'h00);
    
    // -------------------- Data Bus Multiplexer --------------------
    // This always block selects which memory module provides data
    // to the data bus based on the current address.
    
    reg [7:0] mem_data_in;
    
    always @(*) begin
        if (mem_data_from_rom) begin
            // Read from ROM
            mem_data_in = rom_data_out;
        end else if (mem_data_from_ram) begin
            // Read from RAM
            mem_data_in = ram_data_out;
        end else begin
            // No memory selected - high impedance
            mem_data_in = 8'hZZ;
        end
    end
    
    // -------------------- Data Bus Driver --------------------
    // The data bus is bidirectional. It is driven by the CPU
    // when writing to memory, and high-impedance otherwise.
    
    assign data_bus = (mem_write) ? acc_reg : 8'hZZ;
    
    // -------------------- Memory Read Signal --------------------
    // This signal indicates a memory read operation.
    
    assign mem_read = mem_data_from_rom || mem_data_from_ram;
    
    // =========================================================================
    // Output Assignments
    // =========================================================================
    
    assign acc_out = acc_reg;
    assign pc_out = pc_reg;
    assign flags_out = flags_reg;
    assign x_out = x_reg;
    assign y_out = y_reg;
    
    // The CPU runs continuously in this implementation
    assign halt = 1'b0;
    
    // =========================================================================
    // Debug Monitor
    // =========================================================================
    // This always block monitors CPU state and displays information
    // for debugging purposes. It shows register contents when the
    // CPU is reset and on instruction completion.
    
    always @(posedge clk) begin
        if (reset) begin
            // Display initial CPU state on reset
            $display("CPU Reset - PC=%h, ACC=%h, X=%h, Y=%h, FLAGS=%h", 
                     pc_reg, acc_reg, x_reg, y_reg, flags_reg);
        end else begin
            // Display state on instruction completion
            if (done) begin
                $display("PC=%h: opcode=%h, ACC=%h, X=%h, Y=%h, FLAGS=%h",
                         pc_reg, data_bus, acc_reg, x_reg, y_reg, flags_reg);
            end
        end
    end

endmodule
