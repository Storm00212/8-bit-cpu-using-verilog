// ============================================================================
// CPU Testbench - Simple Version
// ============================================================================
// 
// This testbench verifies basic CPU functionality by testing individual
// instructions in sequence without infinite loops.
// ============================================================================

`timescale 1ns/1ps

`include "instructions.vh"

module cpu_tb;
    
    // Testbench signals
    reg clk;
    reg reset;
    wire [7:0] data_bus;
    wire [15:0] addr_bus;
    wire mem_read;
    wire mem_write;
    wire [7:0] acc_out;
    wire [15:0] pc_out;
    wire [7:0] flags_out;
    wire [7:0] x_out;
    wire [7:0] y_out;
    wire halt;
    
    // Memory
    reg [7:0] ram [0:65535];
    reg [7:0] rom [0:65535];
    reg [7:0] mem_data_out;
    
    always @(addr_bus) begin
        if (addr_bus < 16'h0100) begin
            mem_data_out = rom[addr_bus];
        end else begin
            mem_data_out = ram[addr_bus];
        end
    end
    
    always @(posedge clk) begin
        if (mem_write) begin
            ram[addr_bus] <= acc_out;
        end
    end
    
    // Clock
    always #5 clk = ~clk;
    
    // CPU
    cpu_top cpu (
        .clk(clk),
        .reset(reset),
        .data_bus(data_bus),
        .addr_bus(addr_bus),
        .mem_read(mem_read),
        .mem_write(mem_write),
        .acc_out(acc_out),
        .pc_out(pc_out),
        .flags_out(flags_out),
        .x_out(x_out),
        .y_out(y_out),
        .halt(halt)
    );
    
    // Data bus driver
    assign data_bus = (mem_read) ? mem_data_out : 8'hZZ;
    
    integer passed = 0;
    integer failed = 0;
    
    task test_op;
        input [7:0] opcode;
        input [7:0] operand;
        input [7:0] expected;
        input [80:0] name;
        begin
            rom[16'h0000] = opcode;
            rom[16'h0001] = operand;
            rom[16'h0002] = 8'h00;  // NOP to stop
            
            reset = 1;
            @(posedge clk) #1;
            reset = 0;
            
            @(posedge clk) #10;  // Execute opcode
            @(posedge clk) #10;  // Execute operand fetch
            
            if (acc_out == expected) begin
                $display("PASS: %s", name);
                passed = passed + 1;
            end else begin
                $display("FAIL: %s - Expected 0x%02h, Got 0x%02h", name, expected, acc_out);
                failed = failed + 1;
            end
        end
    endtask
    
    initial begin
        clk = 0;
        reset = 0;
        
        $display("========================================");
        $display("8-bit CPU Testbench");
        $display("========================================");
        
        #100;
        
        // Test LDA immediate
        rom[16'h0000] = `OPCODE_LDA_IMM;
        rom[16'h0001] = 8'h55;
        rom[16'h0002] = 8'h00;
        
        reset = 1;
        @(posedge clk) #1;
        reset = 0;
        @(posedge clk) #20;
        
        if (acc_out == 8'h55) begin
            $display("PASS: LDA #immediate");
            passed = passed + 1;
        end else begin
            $display("FAIL: LDA #immediate - Expected 55, Got %h", acc_out);
            failed = failed + 1;
        end
        
        // Test ADD immediate
        rom[16'h0000] = `OPCODE_LDA_IMM;
        rom[16'h0001] = 8'h0A;
        rom[16'h0002] = `OPCODE_ADD_IMM;
        rom[16'h0003] = 8'h05;
        rom[16'h0004] = 8'h00;
        
        @(posedge clk) #20;
        
        if (acc_out == 8'h0F) begin
            $display("PASS: ADD immediate (10 + 5 = 15)");
            passed = passed + 1;
        end else begin
            $display("FAIL: ADD immediate - Expected 0F, Got %h", acc_out);
            failed = failed + 1;
        end
        
        // Test SUB immediate
        rom[16'h0000] = `OPCODE_LDA_IMM;
        rom[16'h0001] = 8'h0A;
        rom[16'h0002] = `OPCODE_SUB_IMM;
        rom[16'h0003] = 8'h03;
        rom[16'h0004] = 8'h00;
        
        @(posedge clk) #20;
        
        if (acc_out == 8'h07) begin
            $display("PASS: SUB immediate (10 - 3 = 7)");
            passed = passed + 1;
        end else begin
            $display("FAIL: SUB immediate - Expected 07, Got %h", acc_out);
            failed = failed + 1;
        end
        
        // Test AND immediate
        rom[16'h0000] = `OPCODE_LDA_IMM;
        rom[16'h0001] = 8'hFF;
        rom[16'h0002] = `OPCODE_AND_IMM;
        rom[16'h0003] = 8'h0F;
        rom[16'h0004] = 8'h00;
        
        @(posedge clk) #20;
        
        if (acc_out == 8'h0F) begin
            $display("PASS: AND immediate (FF & 0F = 0F)");
            passed = passed + 1;
        end else begin
            $display("FAIL: AND immediate - Expected 0F, Got %h", acc_out);
            failed = failed + 1;
        end
        
        // Test OR immediate
        rom[16'h0000] = `OPCODE_LDA_IMM;
        rom[16'h0001] = 8'h0F;
        rom[16'h0002] = `OPCODE_OR_IMM;
        rom[16'h0003] = 8'hF0;
        rom[16'h0004] = 8'h00;
        
        @(posedge clk) #20;
        
        if (acc_out == 8'hFF) begin
            $display("PASS: OR immediate (0F | F0 = FF)");
            passed = passed + 1;
        end else begin
            $display("FAIL: OR immediate - Expected FF, Got %h", acc_out);
            failed = failed + 1;
        end
        
        // Test XOR immediate
        rom[16'h0000] = `OPCODE_LDA_IMM;
        rom[16'h0001] = 8'hFF;
        rom[16'h0002] = `OPCODE_XOR_IMM;
        rom[16'h0003] = 8'hFF;
        rom[16'h0004] = 8'h00;
        
        @(posedge clk) #20;
        
        if (acc_out == 8'h00) begin
            $display("PASS: XOR immediate (FF ^ FF = 00)");
            passed = passed + 1;
        end else begin
            $display("FAIL: XOR immediate - Expected 00, Got %h", acc_out);
            failed = failed + 1;
        end
        
        // Test NOT
        rom[16'h0000] = `OPCODE_LDA_IMM;
        rom[16'h0001] = 8'h00;
        rom[16'h0002] = `OPCODE_NOT;
        rom[16'h0003] = 8'h00;
        
        @(posedge clk) #20;
        
        if (acc_out == 8'hFF) begin
            $display("PASS: NOT (~00 = FF)");
            passed = passed + 1;
        end else begin
            $display("FAIL: NOT - Expected FF, Got %h", acc_out);
            failed = failed + 1;
        end
        
        // Test INC
        rom[16'h0000] = `OPCODE_LDA_IMM;
        rom[16'h0001] = 8'h7F;
        rom[16'h0002] = `OPCODE_INC;
        rom[16'h0003] = 8'h00;
        
        @(posedge clk) #20;
        
        if (acc_out == 8'h80) begin
            $display("PASS: INC (7F + 1 = 80)");
            passed = passed + 1;
        end else begin
            $display("FAIL: INC - Expected 80, Got %h", acc_out);
            failed = failed + 1;
        end
        
        // Test DEC
        rom[16'h0000] = `OPCODE_LDA_IMM;
        rom[16'h0001] = 8'h80;
        rom[16'h0002] = `OPCODE_DEC;
        rom[16'h0003] = 8'h00;
        
        @(posedge clk) #20;
        
        if (acc_out == 8'h7F) begin
            $display("PASS: DEC (80 - 1 = 7F)");
            passed = passed + 1;
        end else begin
            $display("FAIL: DEC - Expected 7F, Got %h", acc_out);
            failed = failed + 1;
        end
        
        // Test LDX
        rom[16'h0000] = `OPCODE_LDX_IMM;
        rom[16'h0001] = 8'hAB;
        rom[16'h0002] = 8'h00;
        
        @(posedge clk) #20;
        
        if (x_out == 8'hAB) begin
            $display("PASS: LDX #immediate");
            passed = passed + 1;
        end else begin
            $display("FAIL: LDX #immediate - Expected AB, Got %h", x_out);
            failed = failed + 1;
        end
        
        // Test LDY
        rom[16'h0000] = `OPCODE_LDY_IMM;
        rom[16'h0001] = 8'hCD;
        rom[16'h0002] = 8'h00;
        
        @(posedge clk) #20;
        
        if (y_out == 8'hCD) begin
            $display("PASS: LDY #immediate");
            passed = passed + 1;
        end else begin
            $display("FAIL: LDY #immediate - Expected CD, Got %h", y_out);
            failed = failed + 1;
        end
        
        // Summary
        $display("");
        $display("========================================");
        $display("Test Summary");
        $display("========================================");
        $display("Passed: %0d", passed);
        $display("Failed: %0d", failed);
        $display("========================================");
        
        #100;
        $finish;
    end
    
    // Timeout
    initial begin
        #5000;
        $display("TIMEOUT");
        $finish;
    end
    
endmodule
